magic
tech scmos
timestamp 1698975745
<< nwell >>
rect -25 10 17 38
<< polysilicon >>
rect -12 28 -10 30
rect 0 28 2 30
rect -12 1 -10 20
rect 0 1 2 20
rect -12 -9 -10 -7
rect 0 -9 2 -7
<< ndiffusion >>
rect -19 -7 -17 1
rect -13 -7 -12 1
rect -10 -7 0 1
rect 2 -7 3 1
rect 7 -7 9 1
<< pdiffusion >>
rect -19 20 -17 28
rect -13 20 -12 28
rect -10 20 -9 28
rect -1 20 0 28
rect 2 20 3 28
rect 7 20 9 28
<< metal1 >>
rect -20 36 10 37
rect -20 32 -17 36
rect -13 32 -6 36
rect -2 32 3 36
rect 7 32 10 36
rect -20 31 10 32
rect -17 28 -13 31
rect 3 28 7 31
rect -7 10 -3 20
rect -7 6 17 10
rect 3 1 7 6
rect -17 -10 -13 -7
rect -19 -11 9 -10
rect -19 -15 -17 -11
rect -13 -15 -7 -11
rect -3 -15 3 -11
rect 7 -15 9 -11
rect -19 -17 9 -15
<< ntransistor >>
rect -12 -7 -10 1
rect 0 -7 2 1
<< ptransistor >>
rect -12 20 -10 28
rect 0 20 2 28
<< polycontact >>
rect -16 4 -12 8
rect 2 13 6 17
<< ndcontact >>
rect -17 -7 -13 1
rect 3 -7 7 1
<< pdcontact >>
rect -17 20 -13 28
rect -9 20 -1 28
rect 3 20 7 28
<< psubstratepcontact >>
rect -17 -15 -13 -11
rect -7 -15 -3 -11
rect 3 -15 7 -11
<< nsubstratencontact >>
rect -17 32 -13 36
rect -6 32 -2 36
rect 3 32 7 36
<< labels >>
rlabel metal1 -7 34 -7 34 5 vdd
rlabel metal1 -11 -13 -11 -13 1 gnd
rlabel polycontact 5 15 5 15 1 inB
rlabel metal1 12 8 12 8 7 out
rlabel polycontact -14 6 -14 6 1 inA
<< end >>
