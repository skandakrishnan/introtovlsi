* SPICE3 file created from ripple.ext - technology: scmos

.option scale=1u

.global Vdd Gnd 

.subckt nand_two out inA inB gnd vdd
M1000 vdd inB out vdd pfet w=8 l=2
+  ad=112 pd=60 as=80 ps=36
M1001 out inB a_n10_n7# Gnd nfet w=8 l=2
+  ad=56 pd=30 as=80 ps=36
M1002 out inA vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_n10_n7# inA gnd Gnd nfet w=8 l=2
+  ad=0 pd=0 as=56 ps=30
C0 inB vdd 4.60fF
C1 vdd inA 3.34fF
C2 gnd Gnd 7.52fF
C3 out Gnd 4.14fF
C4 inB Gnd 3.10fF
C5 inA Gnd 4.36fF
.ends

.subckt or orain orbin orout orvdd orgnd
Xnand_two_0 nand0out orain orain orgnd orvdd nand_two
Xnand_two_2 orout nand1out nand0out orgnd orvdd nand_two
Xnand_two_1 nand1out orbin orbin orgnd orvdd nand_two
C0 orvdd orbin 4.21fF
C1 orain Gnd 13.59fF
C2 orgnd Gnd 28.29fF
C3 nand1out Gnd 7.61fF
C4 orbin Gnd 23.22fF
C5 orout Gnd 2.44fF
C6 nand0out Gnd 17.42fF
.ends

.subckt and anda andb andvout andvdd andgnd
Xnand_two_0 nandout anda andb andgnd andvdd nand_two
Xnand_two_1 andvout nandout nandout andgnd andvdd nand_two
C0 andvdd andb 2.46fF
C1 andvdd nandout 2.06fF
C2 nandout Gnd 7.88fF
C3 andgnd Gnd 29.52fF
C4 andb Gnd 8.66fF
C5 anda Gnd 5.83fF
C6 andvdd Gnd 4.51fF
.ends

.subckt carry carryain carrybin carrycin carryout carryvdd carrygnd
Xor_0 and1out and0out or0out carryvdd carrygnd or
Xor_1 and2out or0out carryout carryvdd carrygnd or
Xand_0 carryain carrycin and0out carryvdd carrygnd and
Xand_1 carrybin carrycin and1out carryvdd carrygnd and
Xand_2 carrybin carryain and2out carryvdd carrygnd and
C0 carrygnd carrybin 2.52fF
C1 carryvdd and0out 2.75fF
C2 carryvdd carryain 10.71fF
C3 or0out carryvdd 3.42fF
C4 carryvdd carrycin 19.54fF
C5 carrybin Gnd 4.64fF
C6 carrygnd Gnd 30.27fF
C7 carrycin Gnd 22.93fF
C8 carryain Gnd 13.21fF
C9 and2out Gnd 15.13fF
C10 or0out Gnd 11.41fF
C11 carryout Gnd 3.76fF
C12 and1out Gnd 11.00fF
C13 and0out Gnd 5.72fF
.ends

.subckt transgate trans_clkp trans_vin trans_clkn trans_vout trans_vdd trans_gnd w_n16_15#
M1000 trans_vout trans_clkn trans_vin Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 trans_vout trans_clkp trans_vin w_n16_15# pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
C0 trans_clkp w_n16_15# 4.53fF
C1 trans_vdd w_n16_15# 11.52fF
C2 trans_gnd Gnd 9.12fF
C3 trans_clkn Gnd 7.46fF
C4 trans_vout Gnd 3.95fF
C5 trans_vin Gnd 4.89fF
C6 trans_clkp Gnd 3.89fF
.ends

.subckt invertor inv_vdd inv_vin inv_vout inv_gnd
M1000 inv_vout inv_vin inv_gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 inv_vout inv_vin inv_vdd inv_vdd pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
C0 inv_vdd inv_vin 2.15fF
C1 inv_gnd Gnd 4.00fF
C2 inv_vout Gnd 3.95fF
C3 inv_vin Gnd 5.97fF
.ends

.subckt xor xora xorb xorvout xorvdd xorgnd
Xtransgate_1 invbout invaout xorb xorvout xorvdd xorgnd xorvdd transgate
Xinvertor_0 xorvdd xorb invbout xorgnd invertor
Xinvertor_1 xorvdd xora invaout xorgnd invertor
Xtransgate_0 xorb xora invbout xorvout xorvdd xorgnd xorvdd transgate
C0 xorvdd invbout 3.02fF
C1 xorb xorvdd 3.47fF
C2 xorvdd xorvout 5.92fF
C3 xorgnd xora 2.16fF
C4 xorb Gnd 42.92fF
C5 xora Gnd 11.23fF
C6 invaout Gnd 6.20fF
C7 xorgnd Gnd 24.44fF
C8 invbout Gnd 16.76fF
C9 xorvdd Gnd 4.89fF
C10 xorvout Gnd 21.02fF
.ends

.subckt sum sumain sumbin sumcin sumvout sumvdd sumgnd
Xxor_0 sumain sumbin xor1out sumvdd sumgnd xor
Xxor_1 xor1out sumcin sumvout sumvdd sumgnd xor
C0 sumcin Gnd 2.44fF
C1 sumvout Gnd 3.29fF
C2 sumbin Gnd 3.20fF
C3 sumain Gnd 3.20fF
C4 sumgnd Gnd 33.56fF
C5 xor1out Gnd 6.61fF
.ends

.subckt fa fa_ain fa_bin fa_cin fa_sout fa_cout fa_vdd fa_gnd
Xcarry_0 fa_ain fa_bin fa_cin fa_cout fa_vdd fa_gnd carry
Xsum_0 fa_bin fa_ain fa_cin fa_sout fa_vdd fa_gnd sum
C0 fa_vdd fa_cin 5.53fF
C1 fa_sout Gnd 4.23fF
C2 fa_ain Gnd 9.59fF
C3 fa_bin Gnd 8.73fF
C4 fa_gnd Gnd 38.49fF
C5 fa_cout Gnd 18.80fF
.ends

.subckt ripple fa_four_vdd fa_four_gnd ri_c0 ri_a0 ri_b0 ri_sout0 ri_a1 ri_b1 ri_sout1
+ ri_a2 ri_b2 ri_sout2 ri_a3 ri_b3 ri_sout3 ri_cout
Xfa_0 ri_a0 ri_b0 ri_c0 ri_sout0 ri_c1 fa_four_vdd fa_four_gnd fa
Xfa_1 ri_a1 ri_b1 ri_c1 ri_sout1 ri_c2 fa_four_vdd fa_four_gnd fa
Xfa_2 ri_a2 ri_b2 ri_c2 ri_sout2 ri_c3 fa_four_vdd fa_four_gnd fa
Xfa_3 ri_a3 ri_b3 ri_c3 ri_sout3 ri_cout fa_four_vdd fa_four_gnd fa
C0 ri_sout3 Gnd 11.98fF
C1 ri_a3 Gnd 5.83fF
C2 ri_b3 Gnd 8.65fF
C3 ri_c3 Gnd 30.46fF
C4 ri_cout Gnd 2.82fF
C5 ri_sout2 Gnd 10.34fF
C6 ri_a2 Gnd 5.45fF
C7 ri_b2 Gnd 6.02fF
C8 ri_c2 Gnd 28.76fF
C9 ri_sout1 Gnd 12.22fF
C10 ri_a1 Gnd 2.07fF
C11 ri_b1 Gnd 3.76fF
C12 ri_c1 Gnd 26.13fF
C13 ri_sout0 Gnd 15.28fF
C14 ri_a0 Gnd 6.02fF
C15 ri_b0 Gnd 7.33fF
C16 fa_four_gnd Gnd 394.89fF
C17 ri_c0 Gnd 5.45fF
C18 fa_four_vdd Gnd 14.95fF
.ends

