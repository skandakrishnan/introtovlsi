magic
tech scmos
timestamp 1698975998
<< nwell >>
rect -6 15 21 43
<< polysilicon >>
rect 4 28 6 30
rect 4 4 6 20
rect 4 -2 6 0
<< ndiffusion >>
rect 3 0 4 4
rect 6 0 7 4
<< pdiffusion >>
rect 3 20 4 28
rect 6 20 7 28
<< metal1 >>
rect -6 40 21 41
rect -6 36 14 40
rect 18 36 21 40
rect -6 34 21 36
rect -1 28 3 34
rect 7 14 11 20
rect -6 10 0 14
rect 7 10 21 14
rect 7 4 11 10
rect -1 -3 3 0
rect -6 -4 21 -3
rect -6 -8 0 -4
rect 4 -8 21 -4
rect -6 -9 21 -8
<< ntransistor >>
rect 4 0 6 4
<< ptransistor >>
rect 4 20 6 28
<< polycontact >>
rect 0 10 4 14
<< ndcontact >>
rect -1 0 3 4
rect 7 0 11 4
<< pdcontact >>
rect -1 20 3 28
rect 7 20 11 28
<< psubstratepcontact >>
rect 0 -8 4 -4
<< nsubstratencontact >>
rect 14 36 18 40
<< end >>
