magic
tech scmos
timestamp 1698986016
<< metal2 >>
rect -17 57 -12 61
rect -8 57 280 61
rect -17 31 280 35
rect -17 13 6 17
rect 10 13 280 17
<< m2contact >>
rect -12 57 -8 61
rect -21 31 -17 35
rect 280 31 284 35
rect 6 13 10 17
use invertor  invertor_0 /home/skanda
timestamp 1698975998
transform 1 0 -11 0 1 21
box -6 -9 21 43
use invertor  invertor_1
timestamp 1698975998
transform 1 0 16 0 1 21
box -6 -9 21 43
use invertor  invertor_2
timestamp 1698975998
transform 1 0 43 0 1 21
box -6 -9 21 43
use invertor  invertor_3
timestamp 1698975998
transform 1 0 70 0 1 21
box -6 -9 21 43
use invertor  invertor_4
timestamp 1698975998
transform 1 0 97 0 1 21
box -6 -9 21 43
use invertor  invertor_5
timestamp 1698975998
transform 1 0 124 0 1 21
box -6 -9 21 43
use invertor  invertor_6
timestamp 1698975998
transform 1 0 151 0 1 21
box -6 -9 21 43
use invertor  invertor_7
timestamp 1698975998
transform 1 0 178 0 1 21
box -6 -9 21 43
use invertor  invertor_8
timestamp 1698975998
transform 1 0 205 0 1 21
box -6 -9 21 43
use invertor  invertor_9
timestamp 1698975998
transform 1 0 232 0 1 21
box -6 -9 21 43
use invertor  invertor_10
timestamp 1698975998
transform 1 0 259 0 1 21
box -6 -9 21 43
<< labels >>
rlabel m2contact -10 59 -10 59 5 vcc
rlabel m2contact 282 33 282 33 7 vout
rlabel m2contact 8 15 8 15 1 gnd
<< end >>
