magic
tech scmos
timestamp 1701981095
<< metal1 >>
rect -1669 753 -1646 754
rect -1669 752 -1468 753
rect 1730 752 1741 754
rect -1669 738 4283 752
rect -1669 400 -1646 738
rect -1588 737 4283 738
rect -1541 603 -1534 737
rect -1181 627 -899 632
rect -704 626 -422 631
rect 1730 603 1741 737
rect -1599 585 -1553 592
rect -1112 583 -1048 592
rect -622 584 -547 591
rect -108 585 12 592
rect 1576 584 1681 591
rect -1600 572 -1552 576
rect -1068 571 -1059 575
rect -570 571 -559 575
rect -49 569 -48 573
rect -44 569 5 573
rect -49 568 5 569
rect 1638 571 1679 575
rect -1601 561 -1560 565
rect -1099 561 -1087 565
rect -601 560 -584 564
rect -99 558 6 564
rect 1355 563 1374 564
rect 1355 559 1369 563
rect 1373 559 1374 563
rect 1638 563 1642 571
rect 2137 560 2152 564
rect 1355 558 1374 559
rect -1597 542 -1537 548
rect -1112 540 -1042 548
rect -605 541 -541 547
rect -106 537 31 547
rect 1639 546 1672 547
rect 1337 542 1352 546
rect 1337 540 1356 542
rect 1643 542 1672 546
rect 1639 541 1672 542
rect 2675 460 2680 737
rect -11 438 137 444
rect 38 419 116 427
rect 565 425 584 427
rect 565 421 580 425
rect 841 425 871 427
rect 845 421 871 425
rect 565 419 584 421
rect 2481 418 2535 427
rect -418 407 -396 411
rect 82 406 103 410
rect 2503 405 2534 409
rect -515 400 -511 401
rect -1679 396 -381 400
rect 59 396 64 400
rect -1669 395 -1646 396
rect -515 242 -511 396
rect 91 395 102 399
rect 565 398 589 399
rect 565 394 585 398
rect 803 394 855 398
rect 2994 394 3009 399
rect 42 376 116 383
rect 557 373 642 382
rect 2510 380 2532 381
rect 2180 376 2203 380
rect 2207 376 2208 380
rect 2514 376 2532 380
rect 2510 375 2532 376
rect 3514 294 3518 737
rect -12 271 113 276
rect 51 254 102 261
rect 561 254 583 258
rect 1684 255 1697 259
rect 3315 252 3397 260
rect -516 234 -511 242
rect -443 240 -408 245
rect 81 241 97 245
rect 3348 239 3385 243
rect -516 230 -411 234
rect 57 230 65 234
rect 563 230 582 234
rect 1490 231 1653 234
rect 3026 231 3072 232
rect 1490 230 1675 231
rect -516 60 -511 230
rect 1649 227 1675 230
rect 3026 227 3068 231
rect 3348 231 3352 239
rect 3849 228 3860 232
rect 46 211 99 217
rect 549 211 1470 218
rect 3001 214 3071 215
rect 3001 210 3066 214
rect 3070 210 3071 214
rect 3349 210 3384 214
rect 3001 209 3071 210
rect 550 187 1717 191
rect 550 165 556 187
rect 69 160 557 165
rect 4205 124 4209 737
rect 4314 124 4580 129
rect 1558 97 1747 101
rect 1618 83 1735 86
rect 1618 79 1671 83
rect 1675 79 1735 83
rect 3823 81 3933 90
rect 4379 82 4455 89
rect 1146 66 1162 70
rect 3865 69 3931 73
rect 4431 69 4455 73
rect -516 59 -496 60
rect 2479 59 2501 61
rect -516 55 1163 59
rect 1627 55 1638 59
rect 1714 55 1729 59
rect 2196 55 2220 59
rect 2483 55 2501 59
rect 3865 57 3870 69
rect 4380 58 4404 62
rect 4907 58 4925 62
rect 1620 36 1742 42
rect 2191 36 2302 42
rect 3830 39 3935 45
rect 4388 39 4460 45
rect 3328 -4 4427 0
<< metal2 >>
rect -1087 648 -44 652
rect -1087 565 -1083 648
rect -49 573 -44 648
rect -49 569 -48 573
rect -49 568 -44 569
rect -584 510 -580 560
rect 1373 559 1638 563
rect 1351 542 1352 546
rect 1356 542 1639 546
rect 1643 542 1645 546
rect 57 510 62 522
rect -584 506 62 510
rect 584 421 841 425
rect 2499 399 2503 405
rect 64 344 68 396
rect 589 394 799 398
rect 803 394 804 398
rect 2198 395 2203 399
rect 2207 395 2504 399
rect 2198 394 2504 395
rect 2207 376 2510 380
rect 538 354 895 358
rect 538 344 542 354
rect 64 340 542 344
rect 583 261 1639 262
rect 583 259 1684 261
rect 583 258 1680 259
rect 587 255 1680 258
rect 587 254 1684 255
rect 582 234 1489 236
rect 586 230 1486 234
rect 65 165 69 230
rect 1621 149 1627 254
rect 3072 227 3348 231
rect 3065 210 3066 214
rect 3070 210 3345 214
rect 1621 144 1675 149
rect 1671 83 1675 144
rect 2224 55 2479 59
rect 1638 -10 1642 55
rect 2553 -10 2557 21
rect 4427 0 4431 69
rect 1638 -14 2559 -10
rect 1638 -15 1642 -14
<< m2contact >>
rect -48 569 -44 573
rect -1087 561 -1083 565
rect -584 560 -580 564
rect 1369 559 1373 563
rect 1638 559 1642 563
rect 1352 542 1356 546
rect 1639 542 1643 546
rect 580 421 584 425
rect 841 421 845 425
rect 2499 405 2503 409
rect 64 396 68 400
rect 585 394 589 398
rect 799 394 803 398
rect 2203 395 2207 399
rect 2203 376 2207 380
rect 2510 376 2514 380
rect 583 254 587 258
rect 1680 255 1684 259
rect 65 230 69 234
rect 582 230 586 234
rect 1486 230 1490 234
rect 3068 227 3072 231
rect 3348 227 3352 231
rect 3066 210 3070 214
rect 3345 210 3349 214
rect 65 160 69 165
rect 1671 79 1675 83
rect 4427 69 4431 73
rect 1638 55 1642 59
rect 2220 55 2224 59
rect 2479 55 2483 59
rect 4427 -4 4431 0
use ff  ff_11
timestamp 1701972462
transform 1 0 3407 0 1 209
box -28 -22 446 90
use ff  ff_9
timestamp 1701972462
transform 1 0 1185 0 1 36
box -28 -22 446 90
use ff  ff_8
timestamp 1701972462
transform 1 0 1753 0 1 36
box -28 -22 446 90
use ff  ff_6
timestamp 1701972462
transform 1 0 120 0 1 211
box -28 -22 446 90
use ff  ff_7
timestamp 1701972462
transform 1 0 -385 0 1 211
box -28 -22 446 90
use ff  ff_10
timestamp 1701972462
transform 1 0 2555 0 1 375
box -28 -22 446 90
use ff  ff_0
timestamp 1701972462
transform 1 0 -535 0 1 541
box -28 -22 446 90
use ff  ff_1
timestamp 1701972462
transform 1 0 -1035 0 1 541
box -28 -22 446 90
use ff  ff_2
timestamp 1701972462
transform 1 0 -1537 0 1 542
box -28 -22 446 90
use ff  ff_3
timestamp 1701972462
transform 1 0 1697 0 1 541
box -28 -22 446 90
use ff  ff_4
timestamp 1701972462
transform 1 0 126 0 1 376
box -28 -22 446 90
use ff  ff_5
timestamp 1701972462
transform 1 0 -383 0 1 377
box -28 -22 446 90
use ripple  ripple_0
timestamp 1701972901
transform 1 0 23 0 1 505
box -24 -509 3847 120
use ff  ff_13
timestamp 1701972462
transform 1 0 4471 0 1 39
box -28 -22 446 90
use ff  ff_12
timestamp 1701972462
transform 1 0 3952 0 1 39
box -28 -22 446 90
<< labels >>
rlabel metal1 -39 560 -39 560 1 ffa0
rlabel metal2 -47 638 -47 638 1 ffc0
rlabel metal2 -43 508 -43 508 1 ffb0
rlabel metal1 -570 573 -570 573 1 in_a0
rlabel metal1 -1068 573 -1068 573 1 in_b0
rlabel metal1 -1600 574 -1600 574 3 in_cin
rlabel metal1 -1599 589 -1599 589 3 vdd
rlabel metal1 -1597 545 -1597 545 3 gnd
rlabel metal1 -1601 563 -1601 563 3 clk
rlabel metal2 1407 561 1407 561 1 ff_ins0
rlabel metal1 2152 562 2152 562 1 out_s0
rlabel metal2 721 396 721 396 1 ff_a1
rlabel metal1 -418 409 -418 409 1 in_b1
rlabel metal2 721 356 721 356 1 ff_b1
rlabel metal2 596 232 596 232 1 ff_a2
rlabel metal1 82 408 82 408 1 in_a1
rlabel metal1 81 243 81 243 1 in_a2
rlabel metal1 380 162 380 162 1 ff_b2
rlabel metal1 -443 243 -443 243 1 in_b2
rlabel metal2 2401 57 2401 57 1 ff_a3
rlabel metal1 1714 57 1714 57 1 in_a3
rlabel metal2 2399 -12 2399 -12 1 ff_b3
rlabel metal1 1146 68 1146 68 1 in_b3
rlabel metal2 2200 396 2200 396 1 ff_ins1
rlabel metal1 3008 396 3008 396 1 out_s1
rlabel metal1 3064 229 3064 229 1 ff_ins2
rlabel metal1 3860 230 3860 230 1 out_s2
rlabel metal1 3874 71 3874 71 1 ff_ins3
rlabel metal1 4404 60 4404 60 1 out_s3
rlabel metal1 4412 -2 4412 -2 1 ff_incout
rlabel metal1 4925 60 4925 60 7 out_cout
<< end >>
