* SPICE3 file created from invertor.ext - technology: scmos

.option scale=1u

.global Vdd Gnd 

.subckt invertor inv_vdd inv_vin inv_vout inv_gnd
M1000 inv_vout inv_vin inv_gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 inv_vout inv_vin inv_vdd inv_vdd pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
C0 inv_vin inv_vdd 2.15fF
C1 inv_gnd Gnd 4.00fF
C2 inv_vout Gnd 3.95fF
C3 inv_vin Gnd 5.97fF
.ends

